** Profile: "SCHEMATIC1-TRANSIENT"  [ D:\redmine_svn\cordia\ADC_01\pcb\sim\FDA-PSpiceFiles\SCHEMATIC1\TRANSIENT.sim ] 

** Creating circuit file "TRANSIENT.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\17.4.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100u 0 1n 
.STEP PARAM Rx LIST 1k 1.1k 
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
